module _8BitCLA (clk, rst, Input_1, Input_2, Carry_In, Carry_Out, Result);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] Input_1;
  input  wire [7:0] Input_2;
  input  wire [0:0] Carry_In;
  output  wire [0:0] Carry_Out;
  output  wire [7:0] Result;

  TC_Splitter8 # (.UUID(64'd1363266575867598353 ^ UUID)) Splitter8_0 (.in(wire_77), .out0(wire_23), .out1(wire_60), .out2(wire_59), .out3(wire_18), .out4(wire_63), .out5(wire_52), .out6(wire_65), .out7(wire_43));
  TC_Splitter8 # (.UUID(64'd4545993000488983991 ^ UUID)) Splitter8_1 (.in(wire_92), .out0(wire_39), .out1(wire_21), .out2(wire_53), .out3(wire_38), .out4(wire_34), .out5(wire_15), .out6(wire_0), .out7(wire_30));
  TC_Maker8 # (.UUID(64'd120906030701661114 ^ UUID)) Maker8_2 (.in0(wire_22), .in1(wire_71), .in2(wire_46), .in3(wire_5), .in4(wire_35), .in5(wire_69), .in6(wire_4), .in7(wire_37), .out(wire_68));
  TC_Xor # (.UUID(64'd877556879023395488 ^ UUID), .BIT_WIDTH(64'd1)) Xor_3 (.in0(wire_18), .in1(wire_38), .out(wire_87));
  TC_Or # (.UUID(64'd1882827039840583370 ^ UUID), .BIT_WIDTH(64'd1)) Or_4 (.in0(wire_18), .in1(wire_38), .out(wire_17));
  TC_And # (.UUID(64'd3698748355134587100 ^ UUID), .BIT_WIDTH(64'd1)) And_5 (.in0(wire_18), .in1(wire_38), .out(wire_72));
  TC_Xor # (.UUID(64'd288130193435245152 ^ UUID), .BIT_WIDTH(64'd1)) Xor_6 (.in0(wire_47), .in1(wire_87), .out(wire_5));
  TC_Xor # (.UUID(64'd1570727524041176803 ^ UUID), .BIT_WIDTH(64'd1)) Xor_7 (.in0(wire_59), .in1(wire_53), .out(wire_78));
  TC_Or # (.UUID(64'd3472114504912624526 ^ UUID), .BIT_WIDTH(64'd1)) Or_8 (.in0(wire_59), .in1(wire_53), .out(wire_14));
  TC_And # (.UUID(64'd468728314573900789 ^ UUID), .BIT_WIDTH(64'd1)) And_9 (.in0(wire_59), .in1(wire_53), .out(wire_6));
  TC_Xor # (.UUID(64'd1462376088986015870 ^ UUID), .BIT_WIDTH(64'd1)) Xor_10 (.in0(wire_24), .in1(wire_78), .out(wire_46));
  TC_Xor # (.UUID(64'd956862460110782301 ^ UUID), .BIT_WIDTH(64'd1)) Xor_11 (.in0(wire_60), .in1(wire_21), .out(wire_89));
  TC_Or # (.UUID(64'd2535926241001393682 ^ UUID), .BIT_WIDTH(64'd1)) Or_12 (.in0(wire_60), .in1(wire_21), .out(wire_7));
  TC_And # (.UUID(64'd774416326559536916 ^ UUID), .BIT_WIDTH(64'd1)) And_13 (.in0(wire_60), .in1(wire_21), .out(wire_32));
  TC_Xor # (.UUID(64'd1983300456363222602 ^ UUID), .BIT_WIDTH(64'd1)) Xor_14 (.in0(wire_25), .in1(wire_89), .out(wire_71));
  TC_Xor # (.UUID(64'd1438790523366153256 ^ UUID), .BIT_WIDTH(64'd1)) Xor_15 (.in0(wire_23), .in1(wire_39), .out(wire_61));
  TC_Or # (.UUID(64'd4057213562886838880 ^ UUID), .BIT_WIDTH(64'd1)) Or_16 (.in0(wire_23), .in1(wire_39), .out(wire_16));
  TC_And # (.UUID(64'd78060819577920021 ^ UUID), .BIT_WIDTH(64'd1)) And_17 (.in0(wire_23), .in1(wire_39), .out(wire_26));
  TC_Xor # (.UUID(64'd4205237116016132319 ^ UUID), .BIT_WIDTH(64'd1)) Xor_18 (.in0(wire_9), .in1(wire_61), .out(wire_22));
  TC_And # (.UUID(64'd684419781690876276 ^ UUID), .BIT_WIDTH(64'd1)) And_19 (.in0(wire_9), .in1(wire_16), .out(wire_85));
  TC_Or # (.UUID(64'd821167505062151053 ^ UUID), .BIT_WIDTH(64'd1)) Or_20 (.in0(wire_85), .in1(wire_26), .out(wire_25));
  TC_And3 # (.UUID(64'd4208425112274370200 ^ UUID), .BIT_WIDTH(64'd1)) And3_21 (.in0(wire_16), .in1(wire_9), .in2(wire_7), .out(wire_67));
  TC_And # (.UUID(64'd2012978552449534576 ^ UUID), .BIT_WIDTH(64'd1)) And_22 (.in0(wire_26), .in1(wire_7), .out(wire_81));
  TC_Or3 # (.UUID(64'd3007133565735341568 ^ UUID), .BIT_WIDTH(64'd1)) Or3_23 (.in0(wire_67), .in1(wire_81), .in2(wire_32), .out(wire_24));
  TC_And3 # (.UUID(64'd3368192791981945267 ^ UUID), .BIT_WIDTH(64'd1)) And3_24 (.in0(wire_26), .in1(wire_7), .in2(wire_14), .out(wire_28));
  TC_And # (.UUID(64'd355435439995505246 ^ UUID), .BIT_WIDTH(64'd1)) And_25 (.in0(wire_32), .in1(wire_14), .out(wire_8));
  TC_Or3 # (.UUID(64'd596009634663818747 ^ UUID), .BIT_WIDTH(64'd1)) Or3_26 (.in0(wire_41), .in1(wire_28), .in2(wire_8), .out(wire_62));
  TC_And3 # (.UUID(64'd3372424111391546524 ^ UUID), .BIT_WIDTH(64'd1)) And3_27 (.in0(wire_16), .in1(wire_9), .in2(wire_14), .out(wire_86));
  TC_And # (.UUID(64'd2323925436359033839 ^ UUID), .BIT_WIDTH(64'd1)) And_28 (.in0(wire_7), .in1(wire_86), .out(wire_41));
  TC_Or # (.UUID(64'd1738434039769324932 ^ UUID), .BIT_WIDTH(64'd1)) Or_29 (.in0(wire_62), .in1(wire_6), .out(wire_47));
  TC_And3 # (.UUID(64'd1100332553591757354 ^ UUID), .BIT_WIDTH(64'd1)) And3_30 (.in0(wire_26), .in1(wire_7), .in2(wire_14), .out(wire_84));
  TC_And # (.UUID(64'd310608575423910205 ^ UUID), .BIT_WIDTH(64'd1)) And_31 (.in0(wire_6), .in1(wire_17), .out(wire_45));
  TC_Or3 # (.UUID(64'd1886779919504794997 ^ UUID), .BIT_WIDTH(64'd1)) Or3_32 (.in0(wire_20), .in1(wire_75), .in2(wire_49), .out(wire_73));
  TC_And3 # (.UUID(64'd319102909416141999 ^ UUID), .BIT_WIDTH(64'd1)) And3_33 (.in0(wire_16), .in1(wire_9), .in2(wire_7), .out(wire_93));
  TC_And # (.UUID(64'd2523575967694043691 ^ UUID), .BIT_WIDTH(64'd1)) And_34 (.in0(wire_93), .in1(wire_66), .out(wire_20));
  TC_Or # (.UUID(64'd2974262406507855886 ^ UUID), .BIT_WIDTH(64'd1)) Or_35 (.in0(wire_73), .in1(wire_2), .out(wire_44));
  TC_And # (.UUID(64'd1096119273580005180 ^ UUID), .BIT_WIDTH(64'd1)) And_36 (.in0(wire_14), .in1(wire_17), .out(wire_66));
  TC_And # (.UUID(64'd2391588055822513363 ^ UUID), .BIT_WIDTH(64'd1)) And_37 (.in0(wire_84), .in1(wire_17), .out(wire_75));
  TC_And3 # (.UUID(64'd3922284266095187218 ^ UUID), .BIT_WIDTH(64'd1)) And3_38 (.in0(wire_32), .in1(wire_14), .in2(wire_17), .out(wire_49));
  TC_Or # (.UUID(64'd1852078784140238612 ^ UUID), .BIT_WIDTH(64'd1)) Or_39 (.in0(wire_45), .in1(wire_72), .out(wire_2));
  TC_Xor # (.UUID(64'd2827999916726412701 ^ UUID), .BIT_WIDTH(64'd1)) Xor_40 (.in0(wire_43), .in1(wire_30), .out(wire_57));
  TC_Or # (.UUID(64'd286671238069865305 ^ UUID), .BIT_WIDTH(64'd1)) Or_41 (.in0(wire_43), .in1(wire_30), .out(wire_42));
  TC_And # (.UUID(64'd2513183520184454505 ^ UUID), .BIT_WIDTH(64'd1)) And_42 (.in0(wire_43), .in1(wire_30), .out(wire_31));
  TC_Xor # (.UUID(64'd1013593826874971108 ^ UUID), .BIT_WIDTH(64'd1)) Xor_43 (.in0(wire_40), .in1(wire_57), .out(wire_37));
  TC_Xor # (.UUID(64'd590289430492175024 ^ UUID), .BIT_WIDTH(64'd1)) Xor_44 (.in0(wire_65), .in1(wire_0), .out(wire_64));
  TC_Or # (.UUID(64'd3570343352336658340 ^ UUID), .BIT_WIDTH(64'd1)) Or_45 (.in0(wire_65), .in1(wire_0), .out(wire_10));
  TC_And # (.UUID(64'd2652958110817944893 ^ UUID), .BIT_WIDTH(64'd1)) And_46 (.in0(wire_65), .in1(wire_0), .out(wire_1));
  TC_Xor # (.UUID(64'd3035472790016061854 ^ UUID), .BIT_WIDTH(64'd1)) Xor_47 (.in0(wire_51), .in1(wire_64), .out(wire_4));
  TC_Xor # (.UUID(64'd4496303562134602464 ^ UUID), .BIT_WIDTH(64'd1)) Xor_48 (.in0(wire_52), .in1(wire_15), .out(wire_33));
  TC_Or # (.UUID(64'd2346657256708143021 ^ UUID), .BIT_WIDTH(64'd1)) Or_49 (.in0(wire_52), .in1(wire_15), .out(wire_11));
  TC_And # (.UUID(64'd1214026557850716623 ^ UUID), .BIT_WIDTH(64'd1)) And_50 (.in0(wire_52), .in1(wire_15), .out(wire_19));
  TC_Xor # (.UUID(64'd3317782970258836405 ^ UUID), .BIT_WIDTH(64'd1)) Xor_51 (.in0(wire_56), .in1(wire_33), .out(wire_69));
  TC_Xor # (.UUID(64'd3247693518523708462 ^ UUID), .BIT_WIDTH(64'd1)) Xor_52 (.in0(wire_63), .in1(wire_34), .out(wire_13));
  TC_Or # (.UUID(64'd611312273798191746 ^ UUID), .BIT_WIDTH(64'd1)) Or_53 (.in0(wire_63), .in1(wire_34), .out(wire_27));
  TC_And # (.UUID(64'd1596644142936516563 ^ UUID), .BIT_WIDTH(64'd1)) And_54 (.in0(wire_63), .in1(wire_34), .out(wire_58));
  TC_Xor # (.UUID(64'd2414713128709665523 ^ UUID), .BIT_WIDTH(64'd1)) Xor_55 (.in0(wire_44), .in1(wire_13), .out(wire_35));
  TC_And # (.UUID(64'd4559076961395440445 ^ UUID), .BIT_WIDTH(64'd1)) And_56 (.in0(wire_44), .in1(wire_27), .out(wire_36));
  TC_Or # (.UUID(64'd127174856192908223 ^ UUID), .BIT_WIDTH(64'd1)) Or_57 (.in0(wire_36), .in1(wire_58), .out(wire_56));
  TC_And3 # (.UUID(64'd3920477358262431492 ^ UUID), .BIT_WIDTH(64'd1)) And3_58 (.in0(wire_27), .in1(wire_44), .in2(wire_11), .out(wire_79));
  TC_And # (.UUID(64'd911945586939329077 ^ UUID), .BIT_WIDTH(64'd1)) And_59 (.in0(wire_58), .in1(wire_11), .out(wire_82));
  TC_Or3 # (.UUID(64'd802909966248645433 ^ UUID), .BIT_WIDTH(64'd1)) Or3_60 (.in0(wire_79), .in1(wire_82), .in2(wire_19), .out(wire_51));
  TC_And3 # (.UUID(64'd2938230722902350805 ^ UUID), .BIT_WIDTH(64'd1)) And3_61 (.in0(wire_58), .in1(wire_11), .in2(wire_10), .out(wire_12));
  TC_And # (.UUID(64'd961943667533104433 ^ UUID), .BIT_WIDTH(64'd1)) And_62 (.in0(wire_19), .in1(wire_10), .out(wire_3));
  TC_Or3 # (.UUID(64'd3438773578756317535 ^ UUID), .BIT_WIDTH(64'd1)) Or3_63 (.in0(wire_80), .in1(wire_12), .in2(wire_3), .out(wire_88));
  TC_And3 # (.UUID(64'd1399067744441062494 ^ UUID), .BIT_WIDTH(64'd1)) And3_64 (.in0(wire_27), .in1(wire_44), .in2(wire_10), .out(wire_70));
  TC_And # (.UUID(64'd3409150753195372814 ^ UUID), .BIT_WIDTH(64'd1)) And_65 (.in0(wire_11), .in1(wire_70), .out(wire_80));
  TC_Or # (.UUID(64'd3360618236216780728 ^ UUID), .BIT_WIDTH(64'd1)) Or_66 (.in0(wire_88), .in1(wire_1), .out(wire_40));
  TC_And3 # (.UUID(64'd914916826925623977 ^ UUID), .BIT_WIDTH(64'd1)) And3_67 (.in0(wire_58), .in1(wire_11), .in2(wire_10), .out(wire_48));
  TC_And # (.UUID(64'd1406432443970789734 ^ UUID), .BIT_WIDTH(64'd1)) And_68 (.in0(wire_1), .in1(wire_42), .out(wire_76));
  TC_Or3 # (.UUID(64'd4427252883269800664 ^ UUID), .BIT_WIDTH(64'd1)) Or3_69 (.in0(wire_55), .in1(wire_29), .in2(wire_54), .out(wire_90));
  TC_And3 # (.UUID(64'd4245796227306515762 ^ UUID), .BIT_WIDTH(64'd1)) And3_70 (.in0(wire_27), .in1(wire_44), .in2(wire_11), .out(wire_91));
  TC_And # (.UUID(64'd3563635374389594120 ^ UUID), .BIT_WIDTH(64'd1)) And_71 (.in0(wire_91), .in1(wire_83), .out(wire_55));
  TC_Or # (.UUID(64'd1042825299522689870 ^ UUID), .BIT_WIDTH(64'd1)) Or_72 (.in0(wire_90), .in1(wire_74), .out(wire_50));
  TC_And # (.UUID(64'd2889755240663231052 ^ UUID), .BIT_WIDTH(64'd1)) And_73 (.in0(wire_10), .in1(wire_42), .out(wire_83));
  TC_And # (.UUID(64'd2630565048805289062 ^ UUID), .BIT_WIDTH(64'd1)) And_74 (.in0(wire_48), .in1(wire_42), .out(wire_29));
  TC_And3 # (.UUID(64'd2738463119282934834 ^ UUID), .BIT_WIDTH(64'd1)) And3_75 (.in0(wire_19), .in1(wire_10), .in2(wire_42), .out(wire_54));
  TC_Or # (.UUID(64'd3012235053845478274 ^ UUID), .BIT_WIDTH(64'd1)) Or_76 (.in0(wire_76), .in1(wire_31), .out(wire_74));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  assign wire_9 = Carry_In;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  assign Carry_Out = wire_50;
  wire [0:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [7:0] wire_68;
  assign Result = wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [0:0] wire_76;
  wire [7:0] wire_77;
  assign wire_77 = Input_1;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [0:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [0:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [0:0] wire_91;
  wire [7:0] wire_92;
  assign wire_92 = Input_2;
  wire [0:0] wire_93;

endmodule
